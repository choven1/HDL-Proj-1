module SelectMode(InputBits, PatternSignal);
  output [119:0] InputBits;
  input [119:0] PatternSignal;

  assign InputBits = PatternSignal;
  
endmodule