
module Memory(GRBSeq,Cycle,Go,clk,reset);
	output reg [119:0] GRBSeq;
	output Cycle;
	input	Go, clk, reset;

	reg [4:0]	S, nS;
	reg [25:0] Count, nCount;
	parameter	BLACKOUT=5'b00000;

	always @(posedge clk)
		if(reset) begin
		    Count <= 0;
			S <= BLACKOUT; end
		else if (Count [25]) begin
			S <= nS;
			Count <= nCount; end
		else begin
			S <= S;
			Count <= nCount; end
			
	always @(reset, Count)
    if(reset || Count [25])
		nCount = 0;
	else
		nCount = Count+1;

	always @(S, Go) begin
		if(S==BLACKOUT)
            nS = (Go ? 5'b00001 : BLACKOUT);
		else
			nS=S+1;
	end
	
	always @(S)
		case(S)
          	5'b00000: GRBSeq = 120'h000000_000000_000000_000000_000000;
			5'b00001: GRBSeq = 120'h0000FF_000000_000000_000000_000000;
			5'b00010: GRBSeq = 120'h00000F_0003FF_000000_000000_000000;
			5'b00011: GRBSeq = 120'h000003_00020F_000FFF_000000_000000;
			5'b00100: GRBSeq = 120'h000000_000103_00070F_003FFF_000000;
			5'b00101: GRBSeq = 120'h000000_000000_000103_00070F_00FFFF;
			5'b00110: GRBSeq = 120'h000000_000000_000000_00FF3F_000F0F;
			5'b00111: GRBSeq = 120'h000000_000000_00FF0F_000F07_000303;
			5'b01000: GRBSeq = 120'h000000_00FF03_000F07_000301_000000;
			5'b01001: GRBSeq = 120'h00FF00_000F02_000301_000000_000000;
			5'b01010: GRBSeq = 120'h000F00_03FF00_000000_000000_000000;
			5'b01011: GRBSeq = 120'h000300_020F00_0FFF00_000000_000000;
			5'b01100: GRBSeq = 120'h000000_010300_070F00_3FFF00_000000;
			5'b01101: GRBSeq = 120'h000000_000000_010300_070F00_FFFF00;
			5'b01110: GRBSeq = 120'h000000_000000_000000_FF3F00_0F0F00;
			5'b01111: GRBSeq = 120'h000000_000000_FF0F00_0F0700_030300;
			5'b10000: GRBSeq = 120'h000000_FF0300_0F0700_030100_000000;
			5'b10001: GRBSeq = 120'hFF0000_0F0200_030100_000000_000000;
			5'b10010: GRBSeq = 120'h0F0000_FF0003_000000_000000_000000;
			5'b10011: GRBSeq = 120'h030000_0F0002_FF000F_000000_000000;
			5'b10100: GRBSeq = 120'h000000_030001_0F0007_FF003F_000000;
			5'b10101: GRBSeq = 120'h000000_000000_030001_0F0007_FF00FF;
			5'b10110: GRBSeq = 120'h000000_000000_000000_3F00FF_0F000F;
			5'b10111: GRBSeq = 120'h000000_000000_0F00FF_07000F_030003;
			5'b11000: GRBSeq = 120'h000000_0300FF_07000F_010003_000000;
			5'b11001: GRBSeq = 120'h0000FF_02000F_010003_000000_000000;
			5'b11010: GRBSeq = 120'h00000F_010003_000000_000000_000000;
			5'b11011: GRBSeq = 120'h000003_000000_000000_000000_000000;
			5'b11100: GRBSeq = 120'h000000_000000_000000_000000_000000;
			5'b11101: GRBSeq = 120'h000000_000000_000000_000000_000000;
			5'b11110: GRBSeq = 120'h000000_000000_000000_000000_000000;
			5'b11111: GRBSeq = 120'h000000_000000_000000_000000_000000;
			default:  GRBSeq = 120'h000000_000000_000000_000000_000000; 
		endcase
		
	assign Cycle = Count[25];
endmodule

